`ifndef MAX_DATA_WIDTH

  `define MAX_DATA_WIDTH 128
  `define SS_MAX 8
  
`endif

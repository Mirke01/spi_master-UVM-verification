PK     ! >RH�q  �   [Content_Types].xml �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���j�0E����Ѷ�J�(��ɢ�eh
�*�8�i�����Ĕ�ĥI6y�{5��7F'+Q9��A�g	X�re������YQ�\hg!c[�l<��N�bBj3�@��G� #b�<X�.�ts��s�����"X�a�`��b�1y���:I Y�X7�^�k%R��l�˥�sHIY�ą��ou(+�v�7MP9$�U��kr�;�4�L�cZr��P}I��I��fnt�T�Pv��-�\Ft��h��$8'�i�%*hfxp���'Qs�����#wFX���b)~�;��;3�Ѡ;C m���?�
s̒:��O[%�����Q�{�O��q$����r#吷x�jǎ�  �� PK     ! ���   N   _rels/.rels �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���j�0@���ѽQ���N/c���[IL��j���<��]�aG��ӓ�zs�Fu��]��U��	��^�[��x ����1x�p����f��#I)ʃ�Y���������*D��i")��c$���qU���~3��1��jH[{�=E����~
f?��3-���޲]�Tꓸ2�j)�,l0/%��b�
���z���ŉ�,	�	�/�|f\Z���?6�!Y�_�o�]A�  �� PK     ! ߵL�
  �   word/_rels/document.xml.rels �(�                                                                                                                                                                                                                                                                 ��MK�0���!�ݦ]u�t/"�U+xͦ�l���U��+��ťx�q�0������v���)Ȓ:����
ފ��ڕ��H�ί�V/�i�KԴ=�Hq��a��$ӠՔ�]<�|���j�k�k��4]�0f@~��RAؔ� �����}U����Yt|�B2ǛQd�P#+8$Id�����U����y�>���숽}�mG�$9��e�ٔ�rN��x2ُ������w\�m7�8FSwsJ|������y���   �� PK     ! V�+��  �     word/document.xml�]is�6��3�5�؝����R��x���]O���N��R$$q�kIJ�;��P�#Łъ=`b�$�����=R���>M���U�g�t;�fa�����w�k��:Ȣ �3z޹�U燋����Y7��IJ�0Y՝�yg\�EWQ�pLӠ:K�̫|X��y���aRe����!��^Q�!�*v='ȦA�Y�ߋQ��`�s��������4Ѓ�h���ۄ���1�&ELJWx���{b�ڢ��Gi����(�mJ�~��6%s?J[�S�}���X�0/Ӡf��HI��fR�f����q׷�&ԗd�8�٣G�ՊBJ�S0�4�hB�%���3)����U{�����k٢����P�ȕ�&�yV��b%���X�xIdz� �i��7+���|J=�sV�	�t��4���~�
 �I�Z�t��5�=I�]���^��`.T Kx��Ƃ���Ɯ�l<����>���$SݦkQ��/�[ޖ��XS�����Z�g�
?���۔���:s=
�Ұ{9��2$�G��6 �����u.��0ȣ[�]��[ep���*�uͷ;�Y�hk~�Xl�l��%�/��mU[��*w�t�0�$�v��Ʃ�W%�*_~���Ta�p��'eH�u�U��9���U;J���eMug}�Y��P��Co�~=��|L۠�cB6.	ڞ�9����/�oz0�*�̆qF���I�x4f�)iE�)��D qz��z�dO@x�!�L͗<ޗ���q���%l��AWc]�;�{$�� ���aI٥�!�{ޛ��R" ���&g�Sk�M�lĪL���׮w?�a�A�����GA��v������TU�)k�g&t�5�H�{D�8�]Pq?�jZ���US�±��5U��(8�:�uw��%4]�z�)���(�e�=��y����79�9.�P����i9D�}O�ި?p��I\�}N²{�����:Oٴ�T�>����C�c�������,��A����U}�F��nت#��	���V��y�X$�:�m�G=��ݞd��Y�( ��d���zL����`�� 
� Է�	 &:��\VPa�S��%T���9Pt�q�R%�egg�4�����uSe,��մ?���(��h�Ee��u�pM�S�J��F���d��x�����_��#���|����O�"��<��=����V�c>���O����d�sx�r}u	.�.X<ʂDĊ@�R�۰NBr@H�|��7�U�/�������kY�ģ<*��c���N�+�"ͫX��	�'�h���,b!�B�L� ]���s����u�0mlɈ��G6Ī�=�4���{;��-�VMF��� ��FD(4˶U:I� �U��"Z��*�^I��s�s�n�a^�A�F�D(�nX.d�e��ТķO���ш�)�S>�>�;�߬�@p~^�}|�ś�c�f�� ���S�r�V�"@kk.1��:4�LbW2��X
Et��=նe0sG���+�C�~�*aOq��9:4{�TW�`�N^i����S��uc����7����u����T���T-��J��>�]��\��SD4!�I�<��B�E���#�K5,',��{CEz�$���*�՗)�C�~�m�mrmUL�V{!Ms]Ւ�"��T��>4fQ{=h� ai/fY�۟�MNm� ������k�����t����,rmB�'6<ͳ�C���1�E���$q9B�tM'���֬N�%��<����'�Lt�gYVO��h���Y�|�>ρ�Fhi Tm����}�p8b�=�xr>�$>�"�,��ɦs���^6���Zu�t�N�/f	�Lh�'!lBۢ���Z2�o��6�"��E�gp�6ME��y$yH�+��%�K
�n��d��H�I���8�T+�Y /�����C�U��MhƚVH,Z!����Z�D++�{X�b[��A��6�\ו־ok74�A�.F�)��m��Nh �FǞEt(��ǂ�!#6����I��F�םSښ}���a�����A��m��%A{y�s�MÃ���pn�h�"��L�ɕc�F�)�U��e� ��{��r� ���S=��ޕ�u�B���i��D���{�R��̇��􋒿Z󱒚]S0�� >�g�8�C�#dΑ�����!y��ȫ�Uh��֓���|]�|�h�Q�C�~kY>3�x`��B�Gk�m�9%4�cA��VuC�e��]��Y��c%>!�ox�<s�^�H%��}ȁD
\�n�ԉ�b�:�9v� aC��e�'-s'��8�bvz�cYē��o����?���y������g?�cķM,��#�MA�F��*��,G0=�qu˕+`��{5bG�F�y�(��؉z� �BO�3(\�wdR��xE��\vAp�[p�Q�S@��
��.S`�-M{^�KZ�yy�iPY¸ �Y��	�^t��i��Td�'��B�3s��VG����I��r��ܣ�V��N :�u�ٖ4Pm*�m�TvĴtd�2�ӊ� �@��iDj�64���,�Rswj�Q%�P�Ty�6��]��u�|K'�+�}���A�<���!�Es������N��.v�4��z�Y�v������۞
ꞩy����.� �Q�Dĳ�oЖZۜ���r۬$��TS�y�Lҵ���`����"[���5͖�ZPt;ء�k	�:ð�'����v��o��3LMS���u��؟F��k�,�������b�͢x��"�b�!Xh}���3wF����'7�=��:ky~���u01��<�D� e�|�m���v]�ˢU�9ц5�T�c�f��Y�p����d�3�jg����پn6��n�G�cּK���_���+4j��2���� ��<]'t�Q:�ADKeC}�����hR7��@�����B�u��Q�-cΔ$��U\���D_rgΘfw�G��k2IiV_�  �� PK     ! �����  P     word/theme/theme1.xml�YKoG�W�w����Ŏ-��Pq�w��f�	�Up�T�*�z(Ro=Tm�@�~��T-��
���z�c���T�����ߏ��/^�3tD��<iy��U���Mw��;��!�p`���&Dz��?��"�R�	�Dn�)�nU*҇e,��$�7�"�
�"�ߘU���z%�4�P�c`{c8�>A}��۞2�2�J��>��5�(6��CNd�	t�Y�9?�CK-�j>^e�b� bj	m��g>9]N��N�����kl^�-� S��n����
~�},�t)c��Z{ʳʆ��;�f�a�K����v��i�(6����N��P6l.����t�-�e��|���z��P�h2Z@�x�) Cή8� ߘ&�U)eWF��e��;\� `��M���d�}�up<kx���N��˅%-I_�T���S1��x�㋧��ɽ''�~9������+8	�TϿ�������Wn�,����~��Te೯���ѳo>������2�Oc"�ur�x�9��x=�~�i�b'	%N��q��*���'��ѱpmb{��^߱>��XQ�j[�=�Y��MW����I�.�e��G.ٝ��v�)��4-mhD,5���$!
�=>"�Av�R˯{�\�B�)jc�tI��l�]�1�e�R�m�f�js�b�K�l$Tf.��Yn���
�N�q���kXE.%'·.D:$��n@�t��Kݫz�3�{l�H��ȅ��9/#w���8u�L����H� E1��ʩ�+D�!8Y�[�X�~umߤ���,A��X�}���1M^֎�~|���o�����\�0�~���n�����=w��}i���o��b�]Vϫ6�Yo5������������C5a�4]Y��A���4�a.��1\}BUt��Ԍ�P�C�R.�`�����T�֜^ �����Ű`cf��|N�i�
[�p:a�����QmQZa�S�y�ބj@X_�k��L4df$�~�L�r�!�H#m��!5�ܦ/y�K��lO!m� ��5���F�4Q�2�EI��\9�Ğ�cЪYoz��i��!
�q
��n@��I��Un�+�y�`wZ֪K�D�B�],���l�D,��_o6��� G7ZM������y�CK�C�%+�i��Ǌ��(8F6�֩
�T�;�䚞�P�3���*��}&����=I����nƅfVR���������?#S�i����3��k��p�my\��CJ#���,�AYh�ӿ6k]�Ѭoe<LA�9D�	
�NE��}���
f��+救3��L��L����ջ���P4�&�#n>h�<w� ԅ���|��y���LPF���R�/�
6O��k�j��� ��\�U����/h�T�lv����>b�%�D<�<�.�l4 ���L�f�I���Q�r�].�3tvq\�s��Ž�����r9\]Y,�J�"cf�:�����1S��G��U�3�� �d��?   �� PK     ! ���.  �     word/settings.xml�VYo�6~/��`蹊u�P�Y$>�,⦈S�%�6I����Rb�l���E^j��o��9���3����>���a^�������qᏼ�҈��
�'�+����?}�g
kj�\e��x[����W�3�.D�9�k!��)7}��S]��`�$'��C?
���҈�WK��>#�J��1��zM
��s����L5�\[�}�)� �ڒJ96��l n��{��1���ap�u�B�/�g*)
�<�.@�;����໽���0������Do)��1h9�`yģ��hRG�?;"E�Imݑ\"�n�WVd�.$�)���A�z6:��D|	M�U��g�T��^��K�F5Տ(_iQ��A<è���j���ֿ��Di�[$Q��\U��7�
���N��=���P�����j�,8bp�W�%��>�%9?���z]�'	�>����dn�/ ����x��V� ������{@^��=�����ti� g�%�TK"�����2�0gd����ʋH��y������A~k��eh�����Zh-�MW�?���C��|au����/�L�a�v�A�A�0��'�$	��{�F�0��I�j'm��̃xq�&�q2?�$�d�O"�(�ǧ�4���$r����d�Y,fm�����,�?�;�&��b�X.	�-�
��\>]�����Ȫ�����t�� �<,+��fxm�t���m5�I)L�//\f�b��uՠ{������y�#\����WΊ��?�j^���S��}�����C�)���ý)㜔P�H������\���KTUM�p�Q���Иh�*ᇓ��7Q�E��~��\��C'���H/v���%N�t����N6p����z��F���=.o:���I�ڢ
Ϛ%�&A�Uo��gؖ�$~�V�d��,h:�զ� j�J�`F�z�P"���el+��X�r.T����n���N���W���B:�W��IV��NM���p��I�vmk;"����)\��3M�F��`>N��U��~-F�h>J� Ƌ ��p�����i~�   �� PK     ! t?9z�   (   customXml/_rels/item1.xml.rels �(�                                                                                                                                                                                                                                                                 �ϱ��0�����ho��P��K)t;J�GILc�Xji߾�+t�(���Q���E]1��h��jP>N~��j����.�����G{��J	����D60��o���,W�0��H9X)c�t��l'�_u����ݓ���|P�=�;6��w�#w	�E�v
���d*���yB1��ߪ��	�k���  �� PK     ! �z�f�   U   ( customXml/itemProps1.xml �$ (�                                  ��Ak�0����{j{^CW�t]�ױA���$���36���vꎻH�'��j�aG�!�$�5�N�ָ^�����I�V�ޡ�a_��6�Z�TL>�9�%�0����c\N�hQ!�mوB��l�8���@2��3QҴ�4���k?�����R�����ƣ׳E��=c%�s�ۋ�^��n�`o�m濔�����AM�'к�P��yE�  �� PK     ! ��%�  �     word/styles.xml�]�r��}OU�ŧ��+�DI�զ,ي]��ޕ�}���5�a в������3mIV�\e� �`f������|['�W��1O�������_�������Ջ�A�a�����=�������e^�',@��\G�UQl^�ъ���'�a�ع��:,����hf_��_o�"��I\�������d}P�rG�5��k���(c�@�i��7y�v��g�M�#����D��8���� hG����ItƴHA	��P}Z'�1` fQ��a�Ƒ����s\���k�m����nS���D ��	D�,���E�c���ln�"�_�O��j��?W<-���e�Gq|##ױ �*����¼x��a�Ε�к'ʋ��x������_��|0�[.eے0�-������zKj���|f/�_I�#�1������7u�M��8�`B���P�&�t���Y�����p[ps���`���w�q�}T�e��<��ׅ�q>P�?����<~x>8S���:~/,��0]��Ǌ��s����v�|�l��6�''�JI�x�-b�boJN>J�D�zWW��)�F��6�ex
F���(����k�m����]�
u��Ch�P:~���@'u�Ӈ:���������±x#��lh�/�q,��Ʊx�"t4�E�h�L8�l*��}bQ{7��9�����{xp�=��p�w7�����p�v�=��z��n��^��Hy���}�GS��r6<9鱌��0:����-
���
QN�>�2��2XƷ�L���g�W���;�G��b�YF�E�[����6���t��hsޒa�tA<|%"IP�	Z��+�$1���a�q���,>��s��� ��6I�G�),��@���
�?3P0��A�3�!2hD#eЈ̠���'ո4�q3hD�f����&.�뫎Q���e�e�ݻ��m���tcj���0o�p�
dU���g�q.��>����vHT�z%�K��8��h�ʹvxD��#r����}�d�@{K��\o�E��*�^N{&[�������WX� Wq���A;,��?�嬤�"�U��oX���V�Q��y���	��Є������7�O~�t��EƵ��.?V��r�7��*�c�+5 �O�����C���Ч$�S�޼X�qЭ ��|x���L3��� ^��k2LS	��l�w��IpzO��WD�!vL2�/���23Nc�9T�����y�-h�>eL_S0"��p�ы�q�N��Ր��w�Ų.D�T7$`��a����"�P��$��_���?�������_&4����M1=H�t����Ug/�0�c�)Tg<��x���O�Ox��&tX��`	H6�<ٮӜ��
���
�����Qx%9���,^������P`T4(0*)�W����/ө��_����� 50*��N�Dgyj`T:S`T:S`T:S`T:���r)�tSL�Js5H��&-�zó0�'�|��ې�@��>e|)�੾�� R֨�Ŷ��"�6'k�ĢlAE4LΉjkՄ�,�׮2Swrx7�SFlœ�,}�ۊ|�Zߖ��|Ռ^e�����W�jf6<hY&���l�Yy?K�����벡�f�٤��Rt�xzظZI4,�{Z�c�[V���IOKx�Ӟ��O�]��:̾�
�K?��"��.�[�%��e�O�T�p��Uɳ��~>c���<v{��Q0�dG��Wv�.��}��̎	��x��'@�W��^��-�u��	��7u��4gA+Τ���F���c�pc��w����W$���B��wl�C�Rvt��3.ZA{\���.�
��D+�U���r��vT�vT�������Q!
�Q!�Q!�Q�������Q!���B��B��B��B��B��:���N�
QЎ
!Ў
!Ў�֋�
�q�
�]��8*DA;*�@;*�@;*�@;*�@;*�@9*0wrT��vT�vT�vT}����B{��B{G�(.�
QЎ
!Ў
!Ў
!Ў
!Ў
!P�
̝��B�B�U�,�pTh�sTh����Q!
�Q!�Q!�Q!�Q!�Q!�Q����B��B��B�.}�S����G���������L�~���]���*[e��/��_��'*��ϓ����zW]�:���e�>utχ.�{!�9S >�k	j*�.��-A�7�Rz��:�]ѷn	��iW�U~Y^�"�#`�fj�#�yW����!��5C8�]��f�+������{��lw})@�c�Ď�%K�U��c�%͎З=;B_�(>�0xb�Ph��PnTC7�R��v,���j �N5�r�B�Q#�j����=8���0�TC(g�!��p*�R�TC,՞�Ɲj�L5�r�.�TC,�K5Dp���S����PnT�,M5D�R�TC'��;�ʙj�E���4�F1\3�-�j��	�f��5C�l�f�-��%�U�9.[��fG�˞�/�v�V<�v(4�v(7�q�R��jG�R�˖�T㲥N�q�R'ոl�N5.[j��-�Q���NT㲥N�q�R'ոl�N5.[j��-�Q�˖ڨ����0�T㲥N�qْ�j\��F5.[j��-�Q�˖�T㲥N�q�R'ոl�N5.[j��-�Q�˖ڨ�eKV�q�R'ոl��j\��A�����^�Y�=/�m�����ᄟӌ�<����Gw�wV�c�7̉�����{����P���b�n)i,[��x�ͪ������"6��g�ˡ�摁<Ј�aͩ�8p��*u�y(���/ЬT>�e���^�rfzo���7Ʒ��r�.�/�m>��m���8e��V��l.��{u+�ykY��e�ݗ�;��^r����_�];�0�t�.���pr��M�o��aY�Nn�ؽ.�.]�k2;�:S�R?V�.z����,�@@W�z���Ĥ�k������\�5�J��i�{H���YmZS�b+��S��t2�7HB��$�[lc37�a��y�mb��҃Fl�g)6�OPlo&���v��U����gClj��ئV����h�6�!�j���ڳ�K���W����jN�����E��Tnt@j�ڮ���6O�闒�I��Fj��Bj�����f��t��h=�����l'+cR+{�#��Uj&��Hm�,�V��Ӗ����tX͔�h���ک!�2��H��*5S롑�ɳ�Z�byj���t:���;��<esj��I+hds�,d�<�	��w�3u�FL*�eq�Y�e���ٳW��?��~�;,�H0F�Y��*�y'��R�\������"�R��`ow!O t�Y� �,?�sV���k1O�Bćw�T띩V�.��J�dI�!Կ��O��>'�����{���m$V�L���5��v�D��4��SY����L�p���|G����m.��Z�`�}�z�~+��`TAl/*���-�[�=������T��m���(5����G,q#)��h�"JM�#S���d$���k�tJD�)!�]�>M��f5ɷ.���>&��������%U$ߺ�i�{Fķ�Wϖ�G�k"��%H�'D|������/."��u@w�Dܙ��3��+|H�u1���Æ�g��w)��Wg/Cu�& )2����S��lL�Um��*��2�S�of�E�1-����tt��,����E}(�6�'Dou���6
�r��ʨ��<�����ˍ��01�Yic�G�C5E��*����c��F�+�[%��k��+��V�+���A>��5B�vP��3N�����v�?�	�w��=�?���|�1�6~}=��;�O�i�C]l����ތK8bc����e��ڭ�#�;����5�Z�t�^Zpsy�������fS�C\rZ����9y2�zA�~��e��6
,�M�5 �:q,O�ʇ�ڻ�g�N�0�wVo=��>S�BꚯƦÎ�(/����?b�:�]�?�\�#�j��p��w.���u�}g�o��~�Ha�,�.��+�(dV?\���s�j�*S�h2�&Ru1��*����_����n?��x��|�!�����a���N�u����mm-+���Go(�폞�����&N�2%u&#:�8�g��TY��-�w{��+��Sr�P��Ī�[4V��w�&.c�U�D�L��4��d�/�T�b�s%���r:��/X�����{�o��M��\^u�ǅǠ���W�kO��Fsv�h]W�7�^��G���G����yy%�H�	)�3 ��q��i����  �� PK     ! cWr*�     docProps/core.xml �(�                                                                                                                                                                                                                                                                 ��QO�0��M�M��at����(�$�D�[m(lm���n�!��ķ���&�m��+���v+�$S\�y�M�A#��4Szx��ˋ��)�Fi0N�E�$m�t/��1!�- ���	�3er�|h�DS��s Qޒ��QR
��^�Y��k�U�d��t��[mrd�ܞ-�2?�\�����!��[+�(�VѩP��|���կB��b�ӄ��	�A���џ��k	�՟�����IG����-W
]��h�2F�)��UՁ,w��]���wy��eFh�7[�v����n�W=�v]���t؈��QE4a�_D�,p���>d�;����Q��}�M�nu�0�,�=�?
�}�6��Nq�  �� PK     ! ܡ��   6   ( customXml/item1.xml �$ (�                                  ���N�0�_%�	4���N������K��m�ĮuoO�'�h��>�w�_�W��cj`S���,����/����g��a��}��%ZL*㔪��Yd��Nv�`R�Rލ��<�I�8:�Ol/I��,w�w�w<E��W�����C�Vp�������C�V��'���&8�w��ns_��g�;|4!9���/;hk�W��  �� PK     ! 7�wJ  �     word/fontTable.xmlĔ�n�0��'�,ߗ8?�-j��n������v�Hy�;V1�F�:"�������w�Ϻ";�@YS�x�(�Fؕ2��xZ\�P7+^Y#��@�?ܵ�Қ�70Ѣ����'Qb#5�����di��~�u��������5o�RU��G	c9�1�5[�J��Vl�4M9Y!�ب��5�ֺU� �g]u<͕9b����plٌp3��
��,���$g�\��0F�3"��0������ϔh1��6��e�$TCpw$�}�'���Aډ�{�y��N�D͍cnǫ���-�[�d,�-�|G����tY.�V���Vt�Z5bs��S~�]
�[X��~a�%�łv���Ff�c$�s�_�G�c�����G7Jα�u�L�pY��X�:��;{�c��&K�<ܾ��9�X���+"��F�V�����&X��"�
H�����w�M<)-�|�-y+���$��F�YI������G�uB�Gn�|w��i�5��wƿ>-�_t��>�+�pG���E��/0�  �� PK     ! �ԍ�'  �     word/webSettings.xml���j1 �{��r׬R�,�B)�^J���쬆f2!�ڧo�j��^B&�|Ʉ�-v��D��+9R�7T[�����rp+'�k��C%��r1����e�H)�d��%�JnR
�Rl6�����͆"�øV���6a�ɮ��i��E1�G&^�P�X�d�>u�*��"y���'��Dk)�!��\�o��?���Bk"15i��9���r���f�~�I?`|L���ӣ�r���391�G�I��|\{�z岔�F��D��e��!�E�	K�w�Z����9j��r�����  �� PK     ! ~i-��  �   docProps/app.xml �(�                                                                                                                                                                                                                                                                 �R]O�0|����s�Aў:T�R?�.��eo��ײ��}��T}�O�3�xvl�z�\��1Y��t��zM��aW�u_N.�*e�r�qW1�W����0f��b	�v��s�"�'�6L{fz�����AP�[�7�'�Y�M����4'a�g�˧�^QC��K��1�����TF���tCy���QV��ʆ᥁[5`��@�<P4�_|1��UT:s��=/�
����*s��Ց�����* �[��8�~�6��u߭g���boQQ�1�m1�tp�����r	A�`OSP�(���e�W�ѓ���g��t��w�ݔ�^u�W�?�<����=o�)�(80���Z�- |姊�\�g���m��D��~���t�ix���q�g�   �� PK-      ! >RH�q  �                   [Content_Types].xmlPK-      ! ���   N               �  _rels/.relsPK-      ! ߵL�
  �               �  word/_rels/document.xml.relsPK-      ! V�+��  �               	  word/document.xmlPK-      ! �����  P                 word/theme/theme1.xmlPK-      ! ���.  �               4  word/settings.xmlPK-      ! t?9z�   (               �  customXml/_rels/item1.xml.relsPK-      ! �z�f�   U               �!  customXml/itemProps1.xmlPK-      ! ��%�  �               �"  word/styles.xmlPK-      ! cWr*�                 �3  docProps/core.xmlPK-      ! ܡ��   6               f6  customXml/item1.xmlPK-      ! 7�wJ  �               �7  word/fontTable.xmlPK-      ! �ԍ�'  �               �9  word/webSettings.xmlPK-      ! ~i-��  �               -;  docProps/app.xmlPK      �  �=    
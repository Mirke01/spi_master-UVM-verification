package spi_pkg;

    import uvm_pkg::*;
`include "spi_types.sv"
`include "spi_defines.sv"
`include "uvm_macros.svh"
`include "spi_data_item.sv"
`include "spi_config.sv"
`include "spi_sequencer.sv"
`include "spi_sequence_lib.sv"
`include "spi_slave_driver.sv"
`include "spi_master_driver.sv"
`include "spi_monitor.sv"
`include "spi_agent.sv"
`include "spi_env.sv"


endpackage

typedef enum{
  SINGLE_RD,
  SINGLE_WR,
  BLOCK_RD,
  BLOCK_WR,
  RMW }transaction_type_t;

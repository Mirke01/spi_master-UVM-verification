`include "spi_defines.v"
`include "spi_timescale.v"
`include "spi_errors.v"

module spi_shift (clk, rst, latch, byte_sel, len, lsb, go,
                  pos_edge, neg_edge, rx_negedge, tx_negedge,
                  tip, last, 
                  p_in, p_out, s_clk, s_in, s_out);

  parameter Tp = 1;
  
  input                          clk;          // system clock
  input                          rst;          // reset
  input                    [3:0] latch;        // latch signal for storing the data in shift register
  input                    [3:0] byte_sel;     // byte select signals for storing the data in shift register
  input [`SPI_CHAR_LEN_BITS-1:0] len;          // data len in bits (minus one)
  input                          lsb;          // lbs first on the line
  input                          go;           // start stansfer
  input                          pos_edge;     // recognize posedge of sclk
  input                          neg_edge;     // recognize negedge of sclk
  input                          rx_negedge;   // s_in is sampled on negative edge 
  input                          tx_negedge;   // s_out is driven on negative edge
  output                         tip;          // transfer in progress
  output                         last;         // last bit
  input                   [31:0] p_in;         // parallel in
  output     [`SPI_MAX_CHAR-1:0] p_out;        // parallel out
  input                          s_clk;        // serial clock
  input                          s_in;         // serial in
  output                         s_out;        // serial out
                                               
  reg                            s_out;        
  reg                            tip;
                              
  reg     [`SPI_CHAR_LEN_BITS:0] cnt;          // data bit count
  reg        [`SPI_MAX_CHAR-1:0] data;         // shift register
  wire    [`SPI_CHAR_LEN_BITS:0] tx_bit_pos;   // next bit position
  wire    [`SPI_CHAR_LEN_BITS:0] rx_bit_pos;   // next bit position
  wire                           rx_clk;       // rx clock enable
  //(T.D.)
  //wire                           tx_clk;       // tx clock enable
  reg				 tx_clk;
  
  assign p_out = data;
  
  assign tx_bit_pos = lsb ? {!(|len), len} - cnt : cnt - {{`SPI_CHAR_LEN_BITS{1'b0}},1'b1};
  assign rx_bit_pos = lsb ? {!(|len), len} - (rx_negedge ? cnt + {{`SPI_CHAR_LEN_BITS{1'b0}},1'b1} : cnt) : 
                            (rx_negedge ? cnt : cnt - {{`SPI_CHAR_LEN_BITS{1'b0}},1'b1});
  
  assign last = !(|cnt);
  
  assign rx_clk = (rx_negedge ? neg_edge : pos_edge) && (!last || s_clk);
  //(T.D.)
  //assign tx_clk = (tx_negedge ? neg_edge : pos_edge) && !last;
  always @(tx_negedge or neg_edge or pos_edge or last)
  begin
     `ifdef SPI_MOSI_DELAYED_ERR
         tx_clk = (tx_negedge ? pos_edge : neg_edge) & (!last);
     `else
         tx_clk = (tx_negedge ? neg_edge : pos_edge) && !last;
     `endif
  end
  
  // Character bit counter
  always @(posedge clk or posedge rst)
  begin
    if(rst)
      cnt <= #Tp {`SPI_CHAR_LEN_BITS+1{1'b0}};
    else
      begin
        if(tip)
          cnt <= #Tp pos_edge ? (cnt - {{`SPI_CHAR_LEN_BITS{1'b0}}, 1'b1}) : cnt;
        else
          cnt <= #Tp !(|len) ? {1'b1, {`SPI_CHAR_LEN_BITS{1'b0}}} : {1'b0, len};
      end
  end
  
  // Transfer in progress
  always @(posedge clk or posedge rst)
  begin
    if(rst)
      tip <= #Tp 1'b0;
  else if(go && ~tip)
    tip <= #Tp 1'b1;
  else if(tip && last && pos_edge)
    tip <= #Tp 1'b0;
  end
  
  //(T.D.)
  wire	s_out_enable;
  assign s_out_enable = (tip ? tx_clk : go);
 
  // Sending bits to the line
  always @(posedge clk or posedge rst)
  begin
    if (rst)
      s_out   <= #Tp 1'b0;
    else
      //(T.D.) simplified the loading
      //s_out <= #Tp (tx_clk || !tip) ? data[tx_bit_pos[`SPI_CHAR_LEN_BITS-1:0]] : s_out;
      //if (tx_clk || !tip)
        if (s_out_enable) 
         s_out <= #Tp data[tx_bit_pos[`SPI_CHAR_LEN_BITS-1:0]];
        else
          if (!tip && !go)
            s_out <= #Tp 1'b0;
  end
  
  // Receiving bits from the line
  always @(posedge clk or posedge rst)
  begin
    if (rst)
      data   <= #Tp {`SPI_MAX_CHAR{1'b0}};
`ifdef SPI_MAX_CHAR_128
    `ifdef WRITE_AFTER_GOBSY_ERR
    else if (latch[0] && !tip)
    `else
    else if (latch[0] && !go)
    `endif
    begin
      `ifdef TX0_NO_UPDATE_ERR
      `else
          `ifdef TX0_SWAP_ERR   
             if (byte_sel[3])
                 data[31:24] <= #Tp p_in[23:16];
             if (byte_sel[2])
                 data[23:16] <= #Tp p_in[31:24];
             if (byte_sel[1])
                 data[15:8] <= #Tp p_in[7:0];
             if (byte_sel[0])
                 data[7:0] <= #Tp p_in[15:8];
          `else
             if (byte_sel[3])
                 data[31:24] <= #Tp p_in[31:24];
               if (byte_sel[2])
                 data[23:16] <= #Tp p_in[23:16];
               if (byte_sel[1])
                 data[15:8] <= #Tp p_in[15:8];
               if (byte_sel[0])
                 data[7:0] <= #Tp p_in[7:0];
          `endif
       `endif
    end
    `ifdef WRITE_AFTER_GOBSY_ERR
    else if (latch[1] && !tip)
    `else
    else if (latch[1] && !go)
    `endif
    begin
      `ifdef TX1_NO_UPDATE_ERR
      `else
          `ifdef TX1_SWAP_ERR
             if (byte_sel[3])
                   data[63:56] <= #Tp p_in[23:16];
             if (byte_sel[2])
                   data[55:48] <= #Tp p_in[31:24];
             if (byte_sel[1])
                   data[47:40] <= #Tp p_in[7:0];
             if (byte_sel[0])
                   data[39:32] <= #Tp p_in[15:8];
          `else
             if (byte_sel[3])
                   data[63:56] <= #Tp p_in[31:24];
             if (byte_sel[2])
                   data[55:48] <= #Tp p_in[23:16];
             if (byte_sel[1])
                   data[47:40] <= #Tp p_in[15:8];
             if (byte_sel[0])
                   data[39:32] <= #Tp p_in[7:0];
         `endif
      `endif
    end
    `ifdef WRITE_AFTER_GOBSY_ERR
    else if (latch[2] && !tip)
    `else
    else if (latch[2] && !go)
    `endif
    begin
    `ifdef TX2_NO_UPDATE_ERR
    `else
       `ifdef TX2_SWAP_ERR
            if (byte_sel[3])
                data[95:88] <= #Tp p_in[23:16];
            if (byte_sel[2])
                data[87:80] <= #Tp p_in[31:24];
            if (byte_sel[1])
                data[79:72] <= #Tp p_in[7:0];
            if (byte_sel[0])
                data[71:64] <= #Tp p_in[15:8];
        `else
            if (byte_sel[3])
                data[95:88] <= #Tp p_in[31:24];
            if (byte_sel[2])
                data[87:80] <= #Tp p_in[23:16];
            if (byte_sel[1])
                data[79:72] <= #Tp p_in[15:8];
            if (byte_sel[0])
                data[71:64] <= #Tp p_in[7:0];
        `endif
     `endif
    end
    `ifdef WRITE_AFTER_GOBSY_ERR
    else if (latch[3] && !tip)
    `else
    else if (latch[3] && !go)
    `endif
    begin
      `ifdef TX3_NO_UPDATE_ERR
      `else
          `ifdef TX3_SWAP_ERR
             if (byte_sel[3])
                data[127:120] <= #Tp p_in[23:16];
             if (byte_sel[2])
                data[119:112] <= #Tp p_in[31:24];
             if (byte_sel[1])
                data[111:104] <= #Tp p_in[7:0];
             if (byte_sel[0])
                data[103:96] <= #Tp p_in[15:8];
          `else
             if (byte_sel[3])
                data[127:120] <= #Tp p_in[31:24];
             if (byte_sel[2])
                data[119:112] <= #Tp p_in[23:16];
             if (byte_sel[1])
                data[111:104] <= #Tp p_in[15:8];
             if (byte_sel[0])
                data[103:96] <= #Tp p_in[7:0];
         `endif
      `endif
    end
`else
`ifdef SPI_MAX_CHAR_64
    `ifdef WRITE_AFTER_GOBSY_ERR
    else if (latch[0] && !tip)
    `else
    else if (latch[0] && !go)
    `endif
    begin
      `ifdef TX0_NO_UPDATE_ERR
      `else
         `ifdef TX0_SWAP_ERR
             if (byte_sel[3])
                 data[31:24] <= #Tp p_in[23:16];
             if (byte_sel[2])
                 data[23:16] <= #Tp p_in[31:24];
             if (byte_sel[1])
                 data[15:8] <= #Tp p_in[7:0];
             if (byte_sel[0])
                 data[7:0] <= #Tp p_in[15:8];
         `else
             if (byte_sel[3])
                 data[31:24] <= #Tp p_in[31:24];
             if (byte_sel[2])
                 data[23:16] <= #Tp p_in[23:16];
             if (byte_sel[1])
                 data[15:8] <= #Tp p_in[15:8];
             if (byte_sel[0])
                 data[7:0] <= #Tp p_in[7:0];
         `endif
     `endif
    end
    `ifdef WRITE_AFTER_GOBSY_ERR
    else if (latch[1] && !tip)
    `else
    else if (latch[1] && !go)
    `endif
    begin
      `ifdef TX1_NO_UPDATE_ERR
      `else
         `ifdef TX1_SWAP_ERR
             if (byte_sel[3])
                   data[63:56] <= #Tp p_in[23:16];
             if (byte_sel[2])
                   data[55:48] <= #Tp p_in[31:24];
             if (byte_sel[1])
                   data[47:40] <= #Tp p_in[7:0];
             if (byte_sel[0])
                   data[39:32] <= #Tp p_in[15:8];
          `else
             if (byte_sel[3])
                   data[63:56] <= #Tp p_in[31:24];
             if (byte_sel[2])
                   data[55:48] <= #Tp p_in[23:16];
             if (byte_sel[1])
                   data[47:40] <= #Tp p_in[15:8];
             if (byte_sel[0])
                   data[39:32] <= #Tp p_in[7:0];
         `endif
      `endif
   end
`else
    `ifdef WRITE_AFTER_GOBSY_ERR
    else if (latch[0] && !tip)
    `else
    else if (latch[0] && !go)
    `endif
      begin
      `ifdef TX0_NO_UPDATE_ERR
      `else
         `ifdef TX0_SWAP_ERR
             `ifdef SPI_MAX_CHAR_8
                if (byte_sel[0])
                   data[`SPI_MAX_CHAR-1:0] <= #Tp p_in[`SPI_MAX_CHAR-1:0];
            `endif
            `ifdef SPI_MAX_CHAR_16
                if (byte_sel[0])
                   data[7:0] <= #Tp p_in[`SPI_MAX_CHAR-1:8];
               if (byte_sel[1])
                  data[`SPI_MAX_CHAR-1:8] <= #Tp p_in[7:0];
            `endif
            `ifdef SPI_MAX_CHAR_24
               if (byte_sel[0])
                  data[7:0] <= #Tp p_in[`SPI_MAX_CHAR-1:16];
               if (byte_sel[1])
                  data[15:8] <= #Tp p_in[15:8];
               if (byte_sel[2])
                  data[`SPI_MAX_CHAR-1:16] <= #Tp p_in[7:0];
            `endif
            `ifdef SPI_MAX_CHAR_32
               if (byte_sel[0])
                  data[7:0] <= #Tp p_in[15:8];
               if (byte_sel[1])
                  data[15:8] <= #Tp p_in[7:0];
               if (byte_sel[2])
                  data[23:16] <= #Tp p_in[`SPI_MAX_CHAR-1:24];
               if (byte_sel[3])
                  data[`SPI_MAX_CHAR-1:24] <= #Tp p_in[23:16];
            `endif
         `else // No error in TX0
            `ifdef SPI_MAX_CHAR_8
                if (byte_sel[0])
                   data[`SPI_MAX_CHAR-1:0] <= #Tp p_in[`SPI_MAX_CHAR-1:0];
            `endif
            `ifdef SPI_MAX_CHAR_16
                if (byte_sel[0])
                   data[7:0] <= #Tp p_in[7:0];
               if (byte_sel[1])
                  data[`SPI_MAX_CHAR-1:8] <= #Tp p_in[`SPI_MAX_CHAR-1:8];
            `endif
            `ifdef SPI_MAX_CHAR_24
               if (byte_sel[0])
                  data[7:0] <= #Tp p_in[7:0];
               if (byte_sel[1])
                  data[15:8] <= #Tp p_in[15:8];
               if (byte_sel[2])
                  data[`SPI_MAX_CHAR-1:16] <= #Tp p_in[`SPI_MAX_CHAR-1:16];
            `endif
            `ifdef SPI_MAX_CHAR_32
               if (byte_sel[0])
                  data[7:0] <= #Tp p_in[7:0];
               if (byte_sel[1])
                  data[15:8] <= #Tp p_in[15:8];
               if (byte_sel[2])
                  data[23:16] <= #Tp p_in[23:16];
               if (byte_sel[3])
                  data[`SPI_MAX_CHAR-1:24] <= #Tp p_in[`SPI_MAX_CHAR-1:24];
            `endif
          `endif
      `endif
      end
`endif
`endif
    else
    //(T.D.) simplified the loading
      //data[rx_bit_pos[`SPI_CHAR_LEN_BITS-1:0]] <= #Tp rx_clk ? s_in : data[rx_bit_pos[`SPI_CHAR_LEN_BITS-1:0]];
      if (rx_clk)
      begin
        `ifdef RX_NO_UPDATE_ERR
        `else
           `ifdef RX_SHIFT_ERR
                data[rx_bit_pos[`SPI_CHAR_LEN_BITS-1:0] + 3] <= #Tp s_in;
           `else
	        data[rx_bit_pos[`SPI_CHAR_LEN_BITS-1:0]] <= #Tp s_in;
           `endif
        `endif
      end
  end
  
endmodule


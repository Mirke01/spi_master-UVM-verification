package wb_package;
  import uvm_pkg::*;
  
  `include "wb_define.sv"
  `include "wb_types.sv"
  `include "uvm_macros.svh"
  `include "wb_config.sv"
  `include "wb_seq_item.sv"
  `include "wb_slave_monitor.sv"
  `include "wb_slave_driver.sv"
  `include "wb_slave_sequencer.sv"
  `include "wb_slave_agent.sv"
  `include "wb_master_monitor.sv"
  `include "wb_master_driver.sv"
  `include "wb_master_sequencer.sv"
  `include "wb_master_agent.sv"
  `include "wb_env.sv"
  
endpackage
